module nand_gate(
    input a,
    input b,
    output y
);

    assign y = ~(a & b);

endmodule


// TEST-BENCH //

`timescale 1ns / 1ps

module tb_nand_gate;

    reg a;
    reg b;
    wire y;

    nand_gate uut (
        .a(a),
        .b(b),
        .y(y)
    );

    initial begin
        a = 0; b = 0; #10;
        a = 0; b = 1; #10;
        a = 1; b = 0; #10;
        a = 1; b = 1; #10;
        $stop;
    end

endmodule
